    Mac OS X            	   2         �                                      ATTR       �   �                     �     com.apple.quarantine q/0041;5265c9df;Firefox; 