library IEEE;
use IEEE.std_logic_1164.all;

package array_port is
type array_bit is array(natural range <>) of std_logic;
end array_port;
